library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_unsigned.all;
use work.ReedSolomon_package.all;

entity SymbolPowerDecoder is port( 
    in_pow: in data_bus;
    out_dec: out data_bus);
end entity;

architecture RTL of SymbolPowerDecoder is
begin

    with in_pow select out_dec <= 
        "00000001" when "00000000",
        "00000010" when "00000001",
        "00000100" when "00000010",
        "00001000" when "00000011",
        "00010000" when "00000100",
        "00100000" when "00000101",
        "01000000" when "00000110",
        "10000000" when "00000111",
        "01110001" when "00001000",
        "11100010" when "00001001",
        "10110101" when "00001010",
        "00011011" when "00001011",
        "00110110" when "00001100",
        "01101100" when "00001101",
        "11011000" when "00001110",
        "11000001" when "00001111",
        "11110011" when "00010000",
        "10010111" when "00010001",
        "01011111" when "00010010",
        "10111110" when "00010011",
        "00001101" when "00010100",
        "00011010" when "00010101",
        "00110100" when "00010110",
        "01101000" when "00010111",
        "11010000" when "00011000",
        "11010001" when "00011001",
        "11010011" when "00011010",
        "11010111" when "00011011",
        "11011111" when "00011100",
        "11001111" when "00011101",
        "11101111" when "00011110",
        "10101111" when "00011111",
        "00101111" when "00100000",
        "01011110" when "00100001",
        "10111100" when "00100010",
        "00001001" when "00100011",
        "00010010" when "00100100",
        "00100100" when "00100101",
        "01001000" when "00100110",
        "10010000" when "00100111",
        "01010001" when "00101000",
        "10100010" when "00101001",
        "00110101" when "00101010",
        "01101010" when "00101011",
        "11010100" when "00101100",
        "11011001" when "00101101",
        "11000011" when "00101110",
        "11110111" when "00101111",
        "10011111" when "00110000",
        "01001111" when "00110001",
        "10011110" when "00110010",
        "01001101" when "00110011",
        "10011010" when "00110100",
        "01000101" when "00110101",
        "10001010" when "00110110",
        "01100101" when "00110111",
        "11001010" when "00111000",
        "11100101" when "00111001",
        "10111011" when "00111010",
        "00000111" when "00111011",
        "00001110" when "00111100",
        "00011100" when "00111101",
        "00111000" when "00111110",
        "01110000" when "00111111",
        "11100000" when "01000000",
        "10110001" when "01000001",
        "00010011" when "01000010",
        "00100110" when "01000011",
        "01001100" when "01000100",
        "10011000" when "01000101",
        "01000001" when "01000110",
        "10000010" when "01000111",
        "01110101" when "01001000",
        "11101010" when "01001001",
        "10100101" when "01001010",
        "00111011" when "01001011",
        "01110110" when "01001100",
        "11101100" when "01001101",
        "10101001" when "01001110",
        "00100011" when "01001111",
        "01000110" when "01010000",
        "10001100" when "01010001",
        "01101001" when "01010010",
        "11010010" when "01010011",
        "11010101" when "01010100",
        "11011011" when "01010101",
        "11000111" when "01010110",
        "11111111" when "01010111",
        "10001111" when "01011000",
        "01101111" when "01011001",
        "11011110" when "01011010",
        "11001101" when "01011011",
        "11101011" when "01011100",
        "10100111" when "01011101",
        "00111111" when "01011110",
        "01111110" when "01011111",
        "11111100" when "01100000",
        "10001001" when "01100001",
        "01100011" when "01100010",
        "11000110" when "01100011",
        "11111101" when "01100100",
        "10001011" when "01100101",
        "01100111" when "01100110",
        "11001110" when "01100111",
        "11101101" when "01101000",
        "10101011" when "01101001",
        "00100111" when "01101010",
        "01001110" when "01101011",
        "10011100" when "01101100",
        "01001001" when "01101101",
        "10010010" when "01101110",
        "01010101" when "01101111",
        "10101010" when "01110000",
        "00100101" when "01110001",
        "01001010" when "01110010",
        "10010100" when "01110011",
        "01011001" when "01110100",
        "10110010" when "01110101",
        "00010101" when "01110110",
        "00101010" when "01110111",
        "01010100" when "01111000",
        "10101000" when "01111001",
        "00100001" when "01111010",
        "01000010" when "01111011",
        "10000100" when "01111100",
        "01111001" when "01111101",
        "11110010" when "01111110",
        "10010101" when "01111111",
        "01011011" when "10000000",
        "10110110" when "10000001",
        "00011101" when "10000010",
        "00111010" when "10000011",
        "01110100" when "10000100",
        "11101000" when "10000101",
        "10100001" when "10000110",
        "00110011" when "10000111",
        "01100110" when "10001000",
        "11001100" when "10001001",
        "11101001" when "10001010",
        "10100011" when "10001011",
        "00110111" when "10001100",
        "01101110" when "10001101",
        "11011100" when "10001110",
        "11001001" when "10001111",
        "11100011" when "10010000",
        "10110111" when "10010001",
        "00011111" when "10010010",
        "00111110" when "10010011",
        "01111100" when "10010100",
        "11111000" when "10010101",
        "10000001" when "10010110",
        "01110011" when "10010111",
        "11100110" when "10011000",
        "10111101" when "10011001",
        "00001011" when "10011010",
        "00010110" when "10011011",
        "00101100" when "10011100",
        "01011000" when "10011101",
        "10110000" when "10011110",
        "00010001" when "10011111",
        "00100010" when "10100000",
        "01000100" when "10100001",
        "10001000" when "10100010",
        "01100001" when "10100011",
        "11000010" when "10100100",
        "11110101" when "10100101",
        "10011011" when "10100110",
        "01000111" when "10100111",
        "10001110" when "10101000",
        "01101101" when "10101001",
        "11011010" when "10101010",
        "11000101" when "10101011",
        "11111011" when "10101100",
        "10000111" when "10101101",
        "01111111" when "10101110",
        "11111110" when "10101111",
        "10001101" when "10110000",
        "01101011" when "10110001",
        "11010110" when "10110010",
        "11011101" when "10110011",
        "11001011" when "10110100",
        "11100111" when "10110101",
        "10111111" when "10110110",
        "00001111" when "10110111",
        "00011110" when "10111000",
        "00111100" when "10111001",
        "01111000" when "10111010",
        "11110000" when "10111011",
        "10010001" when "10111100",
        "01010011" when "10111101",
        "10100110" when "10111110",
        "00111101" when "10111111",
        "01111010" when "11000000",
        "11110100" when "11000001",
        "10011001" when "11000010",
        "01000011" when "11000011",
        "10000110" when "11000100",
        "01111101" when "11000101",
        "11111010" when "11000110",
        "10000101" when "11000111",
        "01111011" when "11001000",
        "11110110" when "11001001",
        "10011101" when "11001010",
        "01001011" when "11001011",
        "10010110" when "11001100",
        "01011101" when "11001101",
        "10111010" when "11001110",
        "00000101" when "11001111",
        "00001010" when "11010000",
        "00010100" when "11010001",
        "00101000" when "11010010",
        "01010000" when "11010011",
        "10100000" when "11010100",
        "00110001" when "11010101",
        "01100010" when "11010110",
        "11000100" when "11010111",
        "11111001" when "11011000",
        "10000011" when "11011001",
        "01110111" when "11011010",
        "11101110" when "11011011",
        "10101101" when "11011100",
        "00101011" when "11011101",
        "01010110" when "11011110",
        "10101100" when "11011111",
        "00101001" when "11100000",
        "01010010" when "11100001",
        "10100100" when "11100010",
        "00111001" when "11100011",
        "01110010" when "11100100",
        "11100100" when "11100101",
        "10111001" when "11100110",
        "00000011" when "11100111",
        "00000110" when "11101000",
        "00001100" when "11101001",
        "00011000" when "11101010",
        "00110000" when "11101011",
        "01100000" when "11101100",
        "11000000" when "11101101",
        "11110001" when "11101110",
        "10010011" when "11101111",
        "01010111" when "11110000",
        "10101110" when "11110001",
        "00101101" when "11110010",
        "01011010" when "11110011",
        "10110100" when "11110100",
        "00011001" when "11110101",
        "00110010" when "11110110",
        "01100100" when "11110111",
        "11001000" when "11111000",
        "11100001" when "11111001",
        "10110011" when "11111010",
        "00010111" when "11111011",
        "00101110" when "11111100",
        "01011100" when "11111101",
        "10111000" when "11111110",
        "--------" when others;    
        
end architecture;
