library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_unsigned.all;
use work.ReedSolomon_package.all;

entity RSDecoderTb is
end entity;

architecture SIM of RSDecoderTb is
    signal clk: std_logic := '1';
	 signal symin: data_bus;
	 signal symout: parity_bus;
	 signal rst: std_logic := '1';
	 signal counter: std_logic_vector(7 downto 0) := "00000000";
begin
process (clk) begin
	if(falling_edge(clk)) then
		counter <= counter +1;
	end if;
end process;
	with counter select symin <=
	"00000000" when "00000000",

"00000001" when "00000001",

"00000010" when "00000010",

"00000011" when "00000011",

"00000100" when "00000100",

"00000101" when "00000101",

"00000110" when "00000110",

"00000111" when "00000111",

"00001000" when "00001000",

"00001001" when "00001001",

"00001010" when "00001010",

"00001011" when "00001011",

"00001100" when "00001100",

"00001101" when "00001101",

"00001110" when "00001110",

"00001111" when "00001111",

"00010000" when "00010000",

"00010001" when "00010001",

"00010010" when "00010010",

"00010011" when "00010011",

"00010100" when "00010100",

"00010101" when "00010101",

"00010110" when "00010110",

"00010111" when "00010111",

"00011000" when "00011000",

"00011001" when "00011001",

"00011010" when "00011010",

"00011011" when "00011011",

"00011100" when "00011100",

"00011101" when "00011101",

"00011110" when "00011110",

"00011111" when "00011111",

"00100000" when "00100000",

"00100001" when "00100001",

"00100010" when "00100010",

"00100011" when "00100011",

"00100100" when "00100100",

"00100101" when "00100101",

"00100110" when "00100110",

"00100111" when "00100111",

"00101000" when "00101000",

"00101001" when "00101001",

"00101010" when "00101010",

"00101011" when "00101011",

"00101100" when "00101100",

"00101101" when "00101101",

"00101110" when "00101110",

"00101111" when "00101111",

"00110000" when "00110000",

"00110001" when "00110001",

"00110010" when "00110010",

"00110011" when "00110011",

"00110100" when "00110100",

"00110101" when "00110101",

"00110110" when "00110110",

"00110111" when "00110111",

"00111000" when "00111000",

"00111001" when "00111001",

"00111010" when "00111010",

"00111011" when "00111011",

"00111100" when "00111100",

"00111101" when "00111101",

"00111110" when "00111110",

"00111111" when "00111111",

"01000000" when "01000000",

"01000001" when "01000001",

"01000010" when "01000010",

"01000011" when "01000011",

"01000100" when "01000100",

"01000101" when "01000101",

"01000110" when "01000110",

"01000111" when "01000111",

"01001000" when "01001000",

"01001001" when "01001001",

"01001010" when "01001010",

"01001011" when "01001011",

"01001100" when "01001100",

"01001101" when "01001101",

"01001110" when "01001110",

"01001111" when "01001111",

"01010000" when "01010000",

"01010001" when "01010001",

"01010010" when "01010010",

"01010011" when "01010011",

"01010100" when "01010100",

"01010101" when "01010101",

"01010110" when "01010110",

"01010111" when "01010111",

"01011000" when "01011000",

"01011001" when "01011001",

"01011010" when "01011010",

"01011011" when "01011011",

"01011100" when "01011100",

"01011101" when "01011101",

"01011110" when "01011110",

"01011111" when "01011111",

"01100000" when "01100000",

"01100001" when "01100001",

"01100010" when "01100010",

"01100011" when "01100011",

"01100100" when "01100100",

"01100101" when "01100101",

"01100110" when "01100110",

"01100111" when "01100111",

"01101000" when "01101000",

"01101001" when "01101001",

"01101010" when "01101010",

"01101011" when "01101011",

"01101100" when "01101100",

"01101101" when "01101101",

"01101110" when "01101110",

"01101111" when "01101111",

"01110000" when "01110000",

"01110001" when "01110001",

"01110010" when "01110010",

"01110011" when "01110011",

"01110100" when "01110100",

"01110101" when "01110101",

"01110110" when "01110110",

"01110111" when "01110111",

"01111000" when "01111000",

"01111001" when "01111001",

"01111010" when "01111010",

"01111011" when "01111011",

"01111100" when "01111100",

"01111101" when "01111101",

"01111110" when "01111110",

"01111111" when "01111111",

"10000000" when "10000000",

"10000001" when "10000001",

"10000010" when "10000010",

"10000011" when "10000011",

"10000100" when "10000100",

"10000101" when "10000101",

"10000110" when "10000110",

"10000111" when "10000111",

"10001000" when "10001000",

"10001001" when "10001001",

"10001010" when "10001010",

"10001011" when "10001011",

"10001100" when "10001100",

"10001101" when "10001101",

"10001110" when "10001110",

"10001111" when "10001111",

"10010000" when "10010000",

"10010001" when "10010001",

"10010010" when "10010010",

"10010011" when "10010011",

"10010100" when "10010100",

"10010101" when "10010101",

"10010110" when "10010110",

"10010111" when "10010111",

"10011000" when "10011000",

"10011001" when "10011001",

"10011010" when "10011010",

"10011011" when "10011011",

"10011100" when "10011100",

"10011101" when "10011101",

"10011110" when "10011110",

"10011111" when "10011111",

"10100000" when "10100000",

"10100001" when "10100001",

"10100010" when "10100010",

"10100011" when "10100011",

"10100100" when "10100100",

"10100101" when "10100101",

"10100110" when "10100110",

"10100111" when "10100111",

"10101000" when "10101000",

"10101001" when "10101001",

"10101010" when "10101010",

"10101011" when "10101011",

"10101100" when "10101100",

"10101101" when "10101101",

"10101110" when "10101110",

"10101111" when "10101111",

"10110000" when "10110000",

"10110001" when "10110001",

"10110010" when "10110010",

"10110011" when "10110011",

"10110100" when "10110100",

"10110101" when "10110101",

"10110110" when "10110110",

"10110111" when "10110111",

"10111000" when "10111000",

"10111001" when "10111001",

"10111010" when "10111010",

"10111011" when "10111011",

"10111100" when "10111100",

"10111101" when "10111101",

"10111110" when "10111110",

"10111111" when "10111111",

"11000000" when "11000000",

"11000001" when "11000001",

"11000010" when "11000010",

"11000011" when "11000011",

"11000100" when "11000100",

"11000101" when "11000101",

"11000110" when "11000110",

"11000111" when "11000111",

"11001000" when "11001000",

"11001001" when "11001001",

"11001010" when "11001010",

"11001011" when "11001011",

"11001100" when "11001100",

"11001101" when "11001101",

"11001110" when "11001110",

"11001111" when "11001111",

"11010000" when "11010000",

"11010001" when "11010001",

"11010010" when "11010010",

"11010011" when "11010011",

"11010100" when "11010100",

"11010101" when "11010101",

"11010110" when "11010110",

"11010111" when "11010111",

"11011000" when "11011000",

"11011001" when "11011001",

"11011010" when "11011010",

"11011011" when "11011011",

"11011100" when "11011100",

"11011101" when "11011101",

"11011110" when "11011110",

"01000001" when "11011111",

"10000100" when "11100000",

"00010001" when "11100001",

"10000011" when "11100010",

"10110001" when "11100011",

"00011111" when "11100100",

"11011011" when "11100101",

"01010011" when "11100110",

"01110100" when "11100111",

"00100001" when "11101000",

"10010011" when "11101001",

"10010110" when "11101010",

"10010110" when "11101011",

"11001101" when "11101100",

"10100111" when "11101101",

"00001110" when "11101110",

"00011101" when "11101111",

"10110101" when "11110000",

"11001000" when "11110001",

"01100110" when "11110010",

"10000100" when "11110011",

"10101111" when "11110100",

"00100010" when "11110101",

"00100101" when "11110110",

"01100100" when "11110111",

"10111000" when "11111000",

"10011100" when "11111001",
"11000110" when "11111010",
"00000110" when "11111011",
"10011111" when "11111100",
"00010111" when "11111101",
"00101110" when "11111110",
"00000000" when others;


    clk <= not clk after 500 ns;
	 rst <= '0' after 10ns;
    decoder: entity work.RSDecoder(RTL) port map(
        clk => clk,
		  rst_a => rst,
		  enable => '1',
		  in_bus => symin,
		  out_bus => symout);

end architecture;