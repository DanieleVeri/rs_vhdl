library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_unsigned.all;
use work.ReedSolomon_package.all;

entity SymbolPowerDecoder is port( 
    in_pow: in data_bus;
    out_dec: out data_bus);
end entity;

architecture RTL of SymbolPowerDecoder is
begin

    with in_pow select out_dec <= 
		"00000001" when "00000000",
		"00000010" when "00000001",
		"00000100" when "00000010",
		"00001000" when "00000011",
		"00010000" when "00000100",
		"00100000" when "00000101",
		"01000000" when "00000110",
		"10000000" when "00000111",
		"00011101" when "00001000",
		"00111010" when "00001001",
		"01110100" when "00001010",
		"11101000" when "00001011",
		"11001101" when "00001100",
		"10000111" when "00001101",
		"00010011" when "00001110",
		"00100110" when "00001111",
		"01001100" when "00010000",
		"10011000" when "00010001",
		"00101101" when "00010010",
		"01011010" when "00010011",
		"10110100" when "00010100",
		"01110101" when "00010101",
		"11101010" when "00010110",
		"11001001" when "00010111",
		"10001111" when "00011000",
		"00000011" when "00011001",
		"00000110" when "00011010",
		"00001100" when "00011011",
		"00011000" when "00011100",
		"00110000" when "00011101",
		"01100000" when "00011110",
		"11000000" when "00011111",
		"10011101" when "00100000",
		"00100111" when "00100001",
		"01001110" when "00100010",
		"10011100" when "00100011",
		"00100101" when "00100100",
		"01001010" when "00100101",
		"10010100" when "00100110",
		"00110101" when "00100111",
		"01101010" when "00101000",
		"11010100" when "00101001",
		"10110101" when "00101010",
		"01110111" when "00101011",
		"11101110" when "00101100",
		"11000001" when "00101101",
		"10011111" when "00101110",
		"00100011" when "00101111",
		"01000110" when "00110000",
		"10001100" when "00110001",
		"00000101" when "00110010",
		"00001010" when "00110011",
		"00010100" when "00110100",
		"00101000" when "00110101",
		"01010000" when "00110110",
		"10100000" when "00110111",
		"01011101" when "00111000",
		"10111010" when "00111001",
		"01101001" when "00111010",
		"11010010" when "00111011",
		"10111001" when "00111100",
		"01101111" when "00111101",
		"11011110" when "00111110",
		"10100001" when "00111111",
		"01011111" when "01000000",
		"10111110" when "01000001",
		"01100001" when "01000010",
		"11000010" when "01000011",
		"10011001" when "01000100",
		"00101111" when "01000101",
		"01011110" when "01000110",
		"10111100" when "01000111",
		"01100101" when "01001000",
		"11001010" when "01001001",
		"10001001" when "01001010",
		"00001111" when "01001011",
		"00011110" when "01001100",
		"00111100" when "01001101",
		"01111000" when "01001110",
		"11110000" when "01001111",
		"11111101" when "01010000",
		"11100111" when "01010001",
		"11010011" when "01010010",
		"10111011" when "01010011",
		"01101011" when "01010100",
		"11010110" when "01010101",
		"10110001" when "01010110",
		"01111111" when "01010111",
		"11111110" when "01011000",
		"11100001" when "01011001",
		"11011111" when "01011010",
		"10100011" when "01011011",
		"01011011" when "01011100",
		"10110110" when "01011101",
		"01110001" when "01011110",
		"11100010" when "01011111",
		"11011001" when "01100000",
		"10101111" when "01100001",
		"01000011" when "01100010",
		"10000110" when "01100011",
		"00010001" when "01100100",
		"00100010" when "01100101",
		"01000100" when "01100110",
		"10001000" when "01100111",
		"00001101" when "01101000",
		"00011010" when "01101001",
		"00110100" when "01101010",
		"01101000" when "01101011",
		"11010000" when "01101100",
		"10111101" when "01101101",
		"01100111" when "01101110",
		"11001110" when "01101111",
		"10000001" when "01110000",
		"00011111" when "01110001",
		"00111110" when "01110010",
		"01111100" when "01110011",
		"11111000" when "01110100",
		"11101101" when "01110101",
		"11000111" when "01110110",
		"10010011" when "01110111",
		"00111011" when "01111000",
		"01110110" when "01111001",
		"11101100" when "01111010",
		"11000101" when "01111011",
		"10010111" when "01111100",
		"00110011" when "01111101",
		"01100110" when "01111110",
		"11001100" when "01111111",
		"10000101" when "10000000",
		"00010111" when "10000001",
		"00101110" when "10000010",
		"01011100" when "10000011",
		"10111000" when "10000100",
		"01101101" when "10000101",
		"11011010" when "10000110",
		"10101001" when "10000111",
		"01001111" when "10001000",
		"10011110" when "10001001",
		"00100001" when "10001010",
		"01000010" when "10001011",
		"10000100" when "10001100",
		"00010101" when "10001101",
		"00101010" when "10001110",
		"01010100" when "10001111",
		"10101000" when "10010000",
		"01001101" when "10010001",
		"10011010" when "10010010",
		"00101001" when "10010011",
		"01010010" when "10010100",
		"10100100" when "10010101",
		"01010101" when "10010110",
		"10101010" when "10010111",
		"01001001" when "10011000",
		"10010010" when "10011001",
		"00111001" when "10011010",
		"01110010" when "10011011",
		"11100100" when "10011100",
		"11010101" when "10011101",
		"10110111" when "10011110",
		"01110011" when "10011111",
		"11100110" when "10100000",
		"11010001" when "10100001",
		"10111111" when "10100010",
		"01100011" when "10100011",
		"11000110" when "10100100",
		"10010001" when "10100101",
		"00111111" when "10100110",
		"01111110" when "10100111",
		"11111100" when "10101000",
		"11100101" when "10101001",
		"11010111" when "10101010",
		"10110011" when "10101011",
		"01111011" when "10101100",
		"11110110" when "10101101",
		"11110001" when "10101110",
		"11111111" when "10101111",
		"11100011" when "10110000",
		"11011011" when "10110001",
		"10101011" when "10110010",
		"01001011" when "10110011",
		"10010110" when "10110100",
		"00110001" when "10110101",
		"01100010" when "10110110",
		"11000100" when "10110111",
		"10010101" when "10111000",
		"00110111" when "10111001",
		"01101110" when "10111010",
		"11011100" when "10111011",
		"10100101" when "10111100",
		"01010111" when "10111101",
		"10101110" when "10111110",
		"01000001" when "10111111",
		"10000010" when "11000000",
		"00011001" when "11000001",
		"00110010" when "11000010",
		"01100100" when "11000011",
		"11001000" when "11000100",
		"10001101" when "11000101",
		"00000111" when "11000110",
		"00001110" when "11000111",
		"00011100" when "11001000",
		"00111000" when "11001001",
		"01110000" when "11001010",
		"11100000" when "11001011",
		"11011101" when "11001100",
		"10100111" when "11001101",
		"01010011" when "11001110",
		"10100110" when "11001111",
		"01010001" when "11010000",
		"10100010" when "11010001",
		"01011001" when "11010010",
		"10110010" when "11010011",
		"01111001" when "11010100",
		"11110010" when "11010101",
		"11111001" when "11010110",
		"11101111" when "11010111",
		"11000011" when "11011000",
		"10011011" when "11011001",
		"00101011" when "11011010",
		"01010110" when "11011011",
		"10101100" when "11011100",
		"01000101" when "11011101",
		"10001010" when "11011110",
		"00001001" when "11011111",
		"00010010" when "11100000",
		"00100100" when "11100001",
		"01001000" when "11100010",
		"10010000" when "11100011",
		"00111101" when "11100100",
		"01111010" when "11100101",
		"11110100" when "11100110",
		"11110101" when "11100111",
		"11110111" when "11101000",
		"11110011" when "11101001",
		"11111011" when "11101010",
		"11101011" when "11101011",
		"11001011" when "11101100",
		"10001011" when "11101101",
		"00001011" when "11101110",
		"00010110" when "11101111",
		"00101100" when "11110000",
		"01011000" when "11110001",
		"10110000" when "11110010",
		"01111101" when "11110011",
		"11111010" when "11110100",
		"11101001" when "11110101",
		"11001111" when "11110110",
		"10000011" when "11110111",
		"00011011" when "11111000",
		"00110110" when "11111001",
		"01101100" when "11111010",
		"11011000" when "11111011",
		"10101101" when "11111100",
		"01000111" when "11111101",
		"10001110" when "11111110",
		"00000001" when "11111111",
		(others => '-') when others;

end architecture;
