library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_unsigned.all;
use work.ReedSolomon_package.all;

entity SymbolPowerEncoder is port( 
    in_pow: in data_bus;
    out_enc: out data_bus);
end entity;

architecture RTL of SymbolPowerEncoder is
begin

    with in_pow select out_enc <=
			"00000000" when "00000000",
			"00000000" when "00000001",
			"00000001" when "00000010",
			"00011001" when "00000011",
			"00000010" when "00000100",
			"00110010" when "00000101",
			"00011010" when "00000110",
			"11000110" when "00000111",
			"00000011" when "00001000",
			"11011111" when "00001001",
			"00110011" when "00001010",
			"11101110" when "00001011",
			"00011011" when "00001100",
			"01101000" when "00001101",
			"11000111" when "00001110",
			"01001011" when "00001111",
			"00000100" when "00010000",
			"01100100" when "00010001",
			"11100000" when "00010010",
			"00001110" when "00010011",
			"00110100" when "00010100",
			"10001101" when "00010101",
			"11101111" when "00010110",
			"10000001" when "00010111",
			"00011100" when "00011000",
			"11000001" when "00011001",
			"01101001" when "00011010",
			"11111000" when "00011011",
			"11001000" when "00011100",
			"00001000" when "00011101",
			"01001100" when "00011110",
			"01110001" when "00011111",
			"00000101" when "00100000",
			"10001010" when "00100001",
			"01100101" when "00100010",
			"00101111" when "00100011",
			"11100001" when "00100100",
			"00100100" when "00100101",
			"00001111" when "00100110",
			"00100001" when "00100111",
			"00110101" when "00101000",
			"10010011" when "00101001",
			"10001110" when "00101010",
			"11011010" when "00101011",
			"11110000" when "00101100",
			"00010010" when "00101101",
			"10000010" when "00101110",
			"01000101" when "00101111",
			"00011101" when "00110000",
			"10110101" when "00110001",
			"11000010" when "00110010",
			"01111101" when "00110011",
			"01101010" when "00110100",
			"00100111" when "00110101",
			"11111001" when "00110110",
			"10111001" when "00110111",
			"11001001" when "00111000",
			"10011010" when "00111001",
			"00001001" when "00111010",
			"01111000" when "00111011",
			"01001101" when "00111100",
			"11100100" when "00111101",
			"01110010" when "00111110",
			"10100110" when "00111111",
			"00000110" when "01000000",
			"10111111" when "01000001",
			"10001011" when "01000010",
			"01100010" when "01000011",
			"01100110" when "01000100",
			"11011101" when "01000101",
			"00110000" when "01000110",
			"11111101" when "01000111",
			"11100010" when "01001000",
			"10011000" when "01001001",
			"00100101" when "01001010",
			"10110011" when "01001011",
			"00010000" when "01001100",
			"10010001" when "01001101",
			"00100010" when "01001110",
			"10001000" when "01001111",
			"00110110" when "01010000",
			"11010000" when "01010001",
			"10010100" when "01010010",
			"11001110" when "01010011",
			"10001111" when "01010100",
			"10010110" when "01010101",
			"11011011" when "01010110",
			"10111101" when "01010111",
			"11110001" when "01011000",
			"11010010" when "01011001",
			"00010011" when "01011010",
			"01011100" when "01011011",
			"10000011" when "01011100",
			"00111000" when "01011101",
			"01000110" when "01011110",
			"01000000" when "01011111",
			"00011110" when "01100000",
			"01000010" when "01100001",
			"10110110" when "01100010",
			"10100011" when "01100011",
			"11000011" when "01100100",
			"01001000" when "01100101",
			"01111110" when "01100110",
			"01101110" when "01100111",
			"01101011" when "01101000",
			"00111010" when "01101001",
			"00101000" when "01101010",
			"01010100" when "01101011",
			"11111010" when "01101100",
			"10000101" when "01101101",
			"10111010" when "01101110",
			"00111101" when "01101111",
			"11001010" when "01110000",
			"01011110" when "01110001",
			"10011011" when "01110010",
			"10011111" when "01110011",
			"00001010" when "01110100",
			"00010101" when "01110101",
			"01111001" when "01110110",
			"00101011" when "01110111",
			"01001110" when "01111000",
			"11010100" when "01111001",
			"11100101" when "01111010",
			"10101100" when "01111011",
			"01110011" when "01111100",
			"11110011" when "01111101",
			"10100111" when "01111110",
			"01010111" when "01111111",
			"00000111" when "10000000",
			"01110000" when "10000001",
			"11000000" when "10000010",
			"11110111" when "10000011",
			"10001100" when "10000100",
			"10000000" when "10000101",
			"01100011" when "10000110",
			"00001101" when "10000111",
			"01100111" when "10001000",
			"01001010" when "10001001",
			"11011110" when "10001010",
			"11101101" when "10001011",
			"00110001" when "10001100",
			"11000101" when "10001101",
			"11111110" when "10001110",
			"00011000" when "10001111",
			"11100011" when "10010000",
			"10100101" when "10010001",
			"10011001" when "10010010",
			"01110111" when "10010011",
			"00100110" when "10010100",
			"10111000" when "10010101",
			"10110100" when "10010110",
			"01111100" when "10010111",
			"00010001" when "10011000",
			"01000100" when "10011001",
			"10010010" when "10011010",
			"11011001" when "10011011",
			"00100011" when "10011100",
			"00100000" when "10011101",
			"10001001" when "10011110",
			"00101110" when "10011111",
			"00110111" when "10100000",
			"00111111" when "10100001",
			"11010001" when "10100010",
			"01011011" when "10100011",
			"10010101" when "10100100",
			"10111100" when "10100101",
			"11001111" when "10100110",
			"11001101" when "10100111",
			"10010000" when "10101000",
			"10000111" when "10101001",
			"10010111" when "10101010",
			"10110010" when "10101011",
			"11011100" when "10101100",
			"11111100" when "10101101",
			"10111110" when "10101110",
			"01100001" when "10101111",
			"11110010" when "10110000",
			"01010110" when "10110001",
			"11010011" when "10110010",
			"10101011" when "10110011",
			"00010100" when "10110100",
			"00101010" when "10110101",
			"01011101" when "10110110",
			"10011110" when "10110111",
			"10000100" when "10111000",
			"00111100" when "10111001",
			"00111001" when "10111010",
			"01010011" when "10111011",
			"01000111" when "10111100",
			"01101101" when "10111101",
			"01000001" when "10111110",
			"10100010" when "10111111",
			"00011111" when "11000000",
			"00101101" when "11000001",
			"01000011" when "11000010",
			"11011000" when "11000011",
			"10110111" when "11000100",
			"01111011" when "11000101",
			"10100100" when "11000110",
			"01110110" when "11000111",
			"11000100" when "11001000",
			"00010111" when "11001001",
			"01001001" when "11001010",
			"11101100" when "11001011",
			"01111111" when "11001100",
			"00001100" when "11001101",
			"01101111" when "11001110",
			"11110110" when "11001111",
			"01101100" when "11010000",
			"10100001" when "11010001",
			"00111011" when "11010010",
			"01010010" when "11010011",
			"00101001" when "11010100",
			"10011101" when "11010101",
			"01010101" when "11010110",
			"10101010" when "11010111",
			"11111011" when "11011000",
			"01100000" when "11011001",
			"10000110" when "11011010",
			"10110001" when "11011011",
			"10111011" when "11011100",
			"11001100" when "11011101",
			"00111110" when "11011110",
			"01011010" when "11011111",
			"11001011" when "11100000",
			"01011001" when "11100001",
			"01011111" when "11100010",
			"10110000" when "11100011",
			"10011100" when "11100100",
			"10101001" when "11100101",
			"10100000" when "11100110",
			"01010001" when "11100111",
			"00001011" when "11101000",
			"11110101" when "11101001",
			"00010110" when "11101010",
			"11101011" when "11101011",
			"01111010" when "11101100",
			"01110101" when "11101101",
			"00101100" when "11101110",
			"11010111" when "11101111",
			"01001111" when "11110000",
			"10101110" when "11110001",
			"11010101" when "11110010",
			"11101001" when "11110011",
			"11100110" when "11110100",
			"11100111" when "11110101",
			"10101101" when "11110110",
			"11101000" when "11110111",
			"01110100" when "11111000",
			"11010110" when "11111001",
			"11110100" when "11111010",
			"11101010" when "11111011",
			"10101000" when "11111100",
			"01010000" when "11111101",
			"01011000" when "11111110",
			"10101111" when "11111111",
			(others => '-') when others;
        
end architecture;
