library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_unsigned.all;

entity ReedSolomon is
end ReedSolomon;

architecture RTL of ReedSolomon is
    
begin
    
end RTL;