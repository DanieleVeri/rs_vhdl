library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_unsigned.all;

entity SymbolPowerDecoder is
    port( 
        in_pow: in data_bus;
        out_enc: out data_bus);
end entity;

architecture RTL of SymbolPowerDecoder is
begin
    with in_pow select
        out_enc <= "00000001" when "00000000",
        out_enc <= "00000010" when "00000001",
        out_enc <= "00000100" when "00000010",
        out_enc <= "00001000" when "00000011",
        out_enc <= "00010000" when "00000100",
        out_enc <= "00100000" when "00000101",
        out_enc <= "01000000" when "00000110",
        out_enc <= "10000000" when "00000111",
        out_enc <= "01110001" when "00001000",
        out_enc <= "11100010" when "00001001",
        out_enc <= "10110101" when "00001010",
        out_enc <= "00011011" when "00001011",
        out_enc <= "00110110" when "00001100",
        out_enc <= "01101100" when "00001101",
        out_enc <= "11011000" when "00001110",
        out_enc <= "11000001" when "00001111",
        out_enc <= "11110011" when "00010000",
        out_enc <= "10010111" when "00010001",
        out_enc <= "01011111" when "00010010",
        out_enc <= "10111110" when "00010011",
        out_enc <= "00001101" when "00010100",
        out_enc <= "00011010" when "00010101",
        out_enc <= "00110100" when "00010110",
        out_enc <= "01101000" when "00010111",
        out_enc <= "11010000" when "00011000",
        out_enc <= "11010001" when "00011001",
        out_enc <= "11010011" when "00011010",
        out_enc <= "11010111" when "00011011",
        out_enc <= "11011111" when "00011100",
        out_enc <= "11001111" when "00011101",
        out_enc <= "11101111" when "00011110",
        out_enc <= "10101111" when "00011111",
        out_enc <= "00101111" when "00100000",
        out_enc <= "01011110" when "00100001",
        out_enc <= "10111100" when "00100010",
        out_enc <= "00001001" when "00100011",
        out_enc <= "00010010" when "00100100",
        out_enc <= "00100100" when "00100101",
        out_enc <= "01001000" when "00100110",
        out_enc <= "10010000" when "00100111",
        out_enc <= "01010001" when "00101000",
        out_enc <= "10100010" when "00101001",
        out_enc <= "00110101" when "00101010",
        out_enc <= "01101010" when "00101011",
        out_enc <= "11010100" when "00101100",
        out_enc <= "11011001" when "00101101",
        out_enc <= "11000011" when "00101110",
        out_enc <= "11110111" when "00101111",
        out_enc <= "10011111" when "00110000",
        out_enc <= "01001111" when "00110001",
        out_enc <= "10011110" when "00110010",
        out_enc <= "01001101" when "00110011",
        out_enc <= "10011010" when "00110100",
        out_enc <= "01000101" when "00110101",
        out_enc <= "10001010" when "00110110",
        out_enc <= "01100101" when "00110111",
        out_enc <= "11001010" when "00111000",
        out_enc <= "11100101" when "00111001",
        out_enc <= "10111011" when "00111010",
        out_enc <= "00000111" when "00111011",
        out_enc <= "00001110" when "00111100",
        out_enc <= "00011100" when "00111101",
        out_enc <= "00111000" when "00111110",
        out_enc <= "01110000" when "00111111",
        out_enc <= "11100000" when "01000000",
        out_enc <= "10110001" when "01000001",
        out_enc <= "00010011" when "01000010",
        out_enc <= "00100110" when "01000011",
        out_enc <= "01001100" when "01000100",
        out_enc <= "10011000" when "01000101",
        out_enc <= "01000001" when "01000110",
        out_enc <= "10000010" when "01000111",
        out_enc <= "01110101" when "01001000",
        out_enc <= "11101010" when "01001001",
        out_enc <= "10100101" when "01001010",
        out_enc <= "00111011" when "01001011",
        out_enc <= "01110110" when "01001100",
        out_enc <= "11101100" when "01001101",
        out_enc <= "10101001" when "01001110",
        out_enc <= "00100011" when "01001111",
        out_enc <= "01000110" when "01010000",
        out_enc <= "10001100" when "01010001",
        out_enc <= "01101001" when "01010010",
        out_enc <= "11010010" when "01010011",
        out_enc <= "11010101" when "01010100",
        out_enc <= "11011011" when "01010101",
        out_enc <= "11000111" when "01010110",
        out_enc <= "11111111" when "01010111",
        out_enc <= "10001111" when "01011000",
        out_enc <= "01101111" when "01011001",
        out_enc <= "11011110" when "01011010",
        out_enc <= "11001101" when "01011011",
        out_enc <= "11101011" when "01011100",
        out_enc <= "10100111" when "01011101",
        out_enc <= "00111111" when "01011110",
        out_enc <= "01111110" when "01011111",
        out_enc <= "11111100" when "01100000",
        out_enc <= "10001001" when "01100001",
        out_enc <= "01100011" when "01100010",
        out_enc <= "11000110" when "01100011",
        out_enc <= "11111101" when "01100100",
        out_enc <= "10001011" when "01100101",
        out_enc <= "01100111" when "01100110",
        out_enc <= "11001110" when "01100111",
        out_enc <= "11101101" when "01101000",
        out_enc <= "10101011" when "01101001",
        out_enc <= "00100111" when "01101010",
        out_enc <= "01001110" when "01101011",
        out_enc <= "10011100" when "01101100",
        out_enc <= "01001001" when "01101101",
        out_enc <= "10010010" when "01101110",
        out_enc <= "01010101" when "01101111",
        out_enc <= "10101010" when "01110000",
        out_enc <= "00100101" when "01110001",
        out_enc <= "01001010" when "01110010",
        out_enc <= "10010100" when "01110011",
        out_enc <= "01011001" when "01110100",
        out_enc <= "10110010" when "01110101",
        out_enc <= "00010101" when "01110110",
        out_enc <= "00101010" when "01110111",
        out_enc <= "01010100" when "01111000",
        out_enc <= "10101000" when "01111001",
        out_enc <= "00100001" when "01111010",
        out_enc <= "01000010" when "01111011",
        out_enc <= "10000100" when "01111100",
        out_enc <= "01111001" when "01111101",
        out_enc <= "11110010" when "01111110",
        out_enc <= "10010101" when "01111111",
        out_enc <= "01011011" when "10000000",
        out_enc <= "10110110" when "10000001",
        out_enc <= "00011101" when "10000010",
        out_enc <= "00111010" when "10000011",
        out_enc <= "01110100" when "10000100",
        out_enc <= "11101000" when "10000101",
        out_enc <= "10100001" when "10000110",
        out_enc <= "00110011" when "10000111",
        out_enc <= "01100110" when "10001000",
        out_enc <= "11001100" when "10001001",
        out_enc <= "11101001" when "10001010",
        out_enc <= "10100011" when "10001011",
        out_enc <= "00110111" when "10001100",
        out_enc <= "01101110" when "10001101",
        out_enc <= "11011100" when "10001110",
        out_enc <= "11001001" when "10001111",
        out_enc <= "11100011" when "10010000",
        out_enc <= "10110111" when "10010001",
        out_enc <= "00011111" when "10010010",
        out_enc <= "00111110" when "10010011",
        out_enc <= "01111100" when "10010100",
        out_enc <= "11111000" when "10010101",
        out_enc <= "10000001" when "10010110",
        out_enc <= "01110011" when "10010111",
        out_enc <= "11100110" when "10011000",
        out_enc <= "10111101" when "10011001",
        out_enc <= "00001011" when "10011010",
        out_enc <= "00010110" when "10011011",
        out_enc <= "00101100" when "10011100",
        out_enc <= "01011000" when "10011101",
        out_enc <= "10110000" when "10011110",
        out_enc <= "00010001" when "10011111",
        out_enc <= "00100010" when "10100000",
        out_enc <= "01000100" when "10100001",
        out_enc <= "10001000" when "10100010",
        out_enc <= "01100001" when "10100011",
        out_enc <= "11000010" when "10100100",
        out_enc <= "11110101" when "10100101",
        out_enc <= "10011011" when "10100110",
        out_enc <= "01000111" when "10100111",
        out_enc <= "10001110" when "10101000",
        out_enc <= "01101101" when "10101001",
        out_enc <= "11011010" when "10101010",
        out_enc <= "11000101" when "10101011",
        out_enc <= "11111011" when "10101100",
        out_enc <= "10000111" when "10101101",
        out_enc <= "01111111" when "10101110",
        out_enc <= "11111110" when "10101111",
        out_enc <= "10001101" when "10110000",
        out_enc <= "01101011" when "10110001",
        out_enc <= "11010110" when "10110010",
        out_enc <= "11011101" when "10110011",
        out_enc <= "11001011" when "10110100",
        out_enc <= "11100111" when "10110101",
        out_enc <= "10111111" when "10110110",
        out_enc <= "00001111" when "10110111",
        out_enc <= "00011110" when "10111000",
        out_enc <= "00111100" when "10111001",
        out_enc <= "01111000" when "10111010",
        out_enc <= "11110000" when "10111011",
        out_enc <= "10010001" when "10111100",
        out_enc <= "01010011" when "10111101",
        out_enc <= "10100110" when "10111110",
        out_enc <= "00111101" when "10111111",
        out_enc <= "01111010" when "11000000",
        out_enc <= "11110100" when "11000001",
        out_enc <= "10011001" when "11000010",
        out_enc <= "01000011" when "11000011",
        out_enc <= "10000110" when "11000100",
        out_enc <= "01111101" when "11000101",
        out_enc <= "11111010" when "11000110",
        out_enc <= "10000101" when "11000111",
        out_enc <= "01111011" when "11001000",
        out_enc <= "11110110" when "11001001",
        out_enc <= "10011101" when "11001010",
        out_enc <= "01001011" when "11001011",
        out_enc <= "10010110" when "11001100",
        out_enc <= "01011101" when "11001101",
        out_enc <= "10111010" when "11001110",
        out_enc <= "00000101" when "11001111",
        out_enc <= "00001010" when "11010000",
        out_enc <= "00010100" when "11010001",
        out_enc <= "00101000" when "11010010",
        out_enc <= "01010000" when "11010011",
        out_enc <= "10100000" when "11010100",
        out_enc <= "00110001" when "11010101",
        out_enc <= "01100010" when "11010110",
        out_enc <= "11000100" when "11010111",
        out_enc <= "11111001" when "11011000",
        out_enc <= "10000011" when "11011001",
        out_enc <= "01110111" when "11011010",
        out_enc <= "11101110" when "11011011",
        out_enc <= "10101101" when "11011100",
        out_enc <= "00101011" when "11011101",
        out_enc <= "01010110" when "11011110",
        out_enc <= "10101100" when "11011111",
        out_enc <= "00101001" when "11100000",
        out_enc <= "01010010" when "11100001",
        out_enc <= "10100100" when "11100010",
        out_enc <= "00111001" when "11100011",
        out_enc <= "01110010" when "11100100",
        out_enc <= "11100100" when "11100101",
        out_enc <= "10111001" when "11100110",
        out_enc <= "00000011" when "11100111",
        out_enc <= "00000110" when "11101000",
        out_enc <= "00001100" when "11101001",
        out_enc <= "00011000" when "11101010",
        out_enc <= "00110000" when "11101011",
        out_enc <= "01100000" when "11101100",
        out_enc <= "11000000" when "11101101",
        out_enc <= "11110001" when "11101110",
        out_enc <= "10010011" when "11101111",
        out_enc <= "01010111" when "11110000",
        out_enc <= "10101110" when "11110001",
        out_enc <= "00101101" when "11110010",
        out_enc <= "01011010" when "11110011",
        out_enc <= "10110100" when "11110100",
        out_enc <= "00011001" when "11110101",
        out_enc <= "00110010" when "11110110",
        out_enc <= "01100100" when "11110111",
        out_enc <= "11001000" when "11111000",
        out_enc <= "11100001" when "11111001",
        out_enc <= "10110011" when "11111010",
        out_enc <= "00010111" when "11111011",
        out_enc <= "00101110" when "11111100",
        out_enc <= "01011100" when "11111101",
        out_enc <= "10111000" when "11111110",
        (others => '-') when others;
end architecture;
