  --Example instantiation for system 'HostBridge'
  HostBridge_inst : HostBridge
    port map(
      out_port_from_the_pio_1 => out_port_from_the_pio_1,
      clk_0 => clk_0,
      in_port_to_the_pio_0 => in_port_to_the_pio_0,
      reset_n => reset_n
    );


