library ieee;
use ieee.numeric_std.all;
use ieee.std_logic_1164.all;

package ReedSolomon_package is

   constant N: integer := 255;
   constant K: integer := 223;
   constant M: integer := 8;
   
   subtype data_bus is std_logic_vector(M-1 downto 0);
	
	type parity_bus is array(N-K-1 downto 0) of data_bus;
	
	constant generator_polynomial : parity_bus := (
		"00101101", -- 45 z**0
		"11011000", -- 216 z**1
		"11101111", -- 239 z**2
		"00011000", -- 24 z**3
		"11111101", -- 253 z**4
		"01101000", -- 104 z**5
		"00011011", -- 27 z**6
		"00101000", -- 40 z**7
		"01101011", -- 107 z**8
		"00110010", -- 50 z**9
		"10100011", -- 163 z**10
		"11010010", -- 210 z**11
		"11100011", -- 227 z**12
		"10000110", -- 134 z**13
		"11100000", -- 224 z**14
		"10011110", -- 158 z**15
		"01110111", -- 119 z**16
		"00001101", -- 13 z**17
		"10011110", -- 158 z**18
		"00000001", -- 1 z**19
		"11101110", -- 238 z**20
		"10100100", -- 164 z**21
		"01010010", -- 82 z**22
		"00101011", -- 43 z**23
		"00001111", -- 15 z**24
		"11101000", -- 232 z**25
		"11110110", -- 246 z**26
		"10001110", -- 142 z**27
		"00110010", -- 50 z**28
		"10111101", -- 189 z**29
		"00011101", -- 29 z**30
		"11101000"); -- 232 z**31

end package;