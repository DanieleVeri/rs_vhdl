library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_unsigned.all;
use work.ReedSolomon_package.all;

entity SymbolPowerEncoder is port( 
    in_pow: in data_bus;
    out_enc: out data_bus);
end entity;

architecture RTL of SymbolPowerEncoder is
begin

    with in_pow select out_enc <=
        "00000000" when "00000000",
        "00000000" when "00000001",
        "00000001" when "00000010",
        "11100111" when "00000011",
        "00000010" when "00000100",
        "11001111" when "00000101",
        "11101000" when "00000110",
        "00111011" when "00000111",
        "00000011" when "00001000",
        "00100011" when "00001001",
        "11010000" when "00001010",
        "10011010" when "00001011",
        "11101001" when "00001100",
        "00010100" when "00001101",
        "00111100" when "00001110",
        "10110111" when "00001111",
        "00000100" when "00010000",
        "10011111" when "00010001",
        "00100100" when "00010010",
        "01000010" when "00010011",
        "11010001" when "00010100",
        "01110110" when "00010101",
        "10011011" when "00010110",
        "11111011" when "00010111",
        "11101010" when "00011000",
        "11110101" when "00011001",
        "00010101" when "00011010",
        "00001011" when "00011011",
        "00111101" when "00011100",
        "10000010" when "00011101",
        "10111000" when "00011110",
        "10010010" when "00011111",
        "00000101" when "00100000",
        "01111010" when "00100001",
        "10100000" when "00100010",
        "01001111" when "00100011",
        "00100101" when "00100100",
        "01110001" when "00100101",
        "01000011" when "00100110",
        "01101010" when "00100111",
        "11010010" when "00101000",
        "11100000" when "00101001",
        "01110111" when "00101010",
        "11011101" when "00101011",
        "10011100" when "00101100",
        "11110010" when "00101101",
        "11111100" when "00101110",
        "00100000" when "00101111",
        "11101011" when "00110000",
        "11010101" when "00110001",
        "11110110" when "00110010",
        "10000111" when "00110011",
        "00010110" when "00110100",
        "00101010" when "00110101",
        "00001100" when "00110110",
        "10001100" when "00110111",
        "00111110" when "00111000",
        "11100011" when "00111001",
        "10000011" when "00111010",
        "01001011" when "00111011",
        "10111001" when "00111100",
        "10111111" when "00111101",
        "10010011" when "00111110",
        "01011110" when "00111111",
        "00000110" when "01000000",
        "01000110" when "01000001",
        "01111011" when "01000010",
        "11000011" when "01000011",
        "10100001" when "01000100",
        "00110101" when "01000101",
        "01010000" when "01000110",
        "10100111" when "01000111",
        "00100110" when "01001000",
        "01101101" when "01001001",
        "01110010" when "01001010",
        "11001011" when "01001011",
        "01000100" when "01001100",
        "00110011" when "01001101",
        "01101011" when "01001110",
        "00110001" when "01001111",
        "11010011" when "01010000",
        "00101000" when "01010001",
        "11100001" when "01010010",
        "10111101" when "01010011",
        "01111000" when "01010100",
        "01101111" when "01010101",
        "11011110" when "01010110",
        "11110000" when "01010111",
        "10011101" when "01011000",
        "01110100" when "01011001",
        "11110011" when "01011010",
        "10000000" when "01011011",
        "11111101" when "01011100",
        "11001101" when "01011101",
        "00100001" when "01011110",
        "00010010" when "01011111",
        "11101100" when "01100000",
        "10100011" when "01100001",
        "11010110" when "01100010",
        "01100010" when "01100011",
        "11110111" when "01100100",
        "00110111" when "01100101",
        "10001000" when "01100110",
        "01100110" when "01100111",
        "00010111" when "01101000",
        "01010010" when "01101001",
        "00101011" when "01101010",
        "10110001" when "01101011",
        "00001101" when "01101100",
        "10101001" when "01101101",
        "10001101" when "01101110",
        "01011001" when "01101111",
        "00111111" when "01110000",
        "00001000" when "01110001",
        "11100100" when "01110010",
        "10010111" when "01110011",
        "10000100" when "01110100",
        "01001000" when "01110101",
        "01001100" when "01110110",
        "11011010" when "01110111",
        "10111010" when "01111000",
        "01111101" when "01111001",
        "11000000" when "01111010",
        "11001000" when "01111011",
        "10010100" when "01111100",
        "11000101" when "01111101",
        "01011111" when "01111110",
        "10101110" when "01111111",
        "00000111" when "10000000",
        "10010110" when "10000001",
        "01000111" when "10000010",
        "11011001" when "10000011",
        "01111100" when "10000100",
        "11000111" when "10000101",
        "11000100" when "10000110",
        "10101101" when "10000111",
        "10100010" when "10001000",
        "01100001" when "10001001",
        "00110110" when "10001010",
        "01100101" when "10001011",
        "01010001" when "10001100",
        "10110000" when "10001101",
        "10101000" when "10001110",
        "01011000" when "10001111",
        "00100111" when "10010000",
        "10111100" when "10010001",
        "01101110" when "10010010",
        "11101111" when "10010011",
        "01110011" when "10010100",
        "01111111" when "10010101",
        "11001100" when "10010110",
        "00010001" when "10010111",
        "01000101" when "10011000",
        "11000010" when "10011001",
        "00110100" when "10011010",
        "10100110" when "10011011",
        "01101100" when "10011100",
        "11001010" when "10011101",
        "00110010" when "10011110",
        "00110000" when "10011111",
        "11010100" when "10100000",
        "10000110" when "10100001",
        "00101001" when "10100010",
        "10001011" when "10100011",
        "11100010" when "10100100",
        "01001010" when "10100101",
        "10111110" when "10100110",
        "01011101" when "10100111",
        "01111001" when "10101000",
        "01001110" when "10101001",
        "01110000" when "10101010",
        "01101001" when "10101011",
        "11011111" when "10101100",
        "11011100" when "10101101",
        "11110001" when "10101110",
        "00011111" when "10101111",
        "10011110" when "10110000",
        "01000001" when "10110001",
        "01110101" when "10110010",
        "11111010" when "10110011",
        "11110100" when "10110100",
        "00001010" when "10110101",
        "10000001" when "10110110",
        "10010001" when "10110111",
        "11111110" when "10111000",
        "11100110" when "10111001",
        "11001110" when "10111010",
        "00111010" when "10111011",
        "00100010" when "10111100",
        "10011001" when "10111101",
        "00010011" when "10111110",
        "10110110" when "10111111",
        "11101101" when "11000000",
        "00001111" when "11000001",
        "10100100" when "11000010",
        "00101110" when "11000011",
        "11010111" when "11000100",
        "10101011" when "11000101",
        "01100011" when "11000110",
        "01010110" when "11000111",
        "11111000" when "11001000",
        "10001111" when "11001001",
        "00111000" when "11001010",
        "10110100" when "11001011",
        "10001001" when "11001100",
        "01011011" when "11001101",
        "01100111" when "11001110",
        "00011101" when "11001111",
        "00011000" when "11010000",
        "00011001" when "11010001",
        "01010011" when "11010010",
        "00011010" when "11010011",
        "00101100" when "11010100",
        "01010100" when "11010101",
        "10110010" when "11010110",
        "00011011" when "11010111",
        "00001110" when "11011000",
        "00101101" when "11011001",
        "10101010" when "11011010",
        "01010101" when "11011011",
        "10001110" when "11011100",
        "10110011" when "11011101",
        "01011010" when "11011110",
        "00011100" when "11011111",
        "01000000" when "11100000",
        "11111001" when "11100001",
        "00001001" when "11100010",
        "10010000" when "11100011",
        "11100101" when "11100100",
        "00111001" when "11100101",
        "10011000" when "11100110",
        "10110101" when "11100111",
        "10000101" when "11101000",
        "10001010" when "11101001",
        "01001001" when "11101010",
        "01011100" when "11101011",
        "01001101" when "11101100",
        "01101000" when "11101101",
        "11011011" when "11101110",
        "00011110" when "11101111",
        "10111011" when "11110000",
        "11101110" when "11110001",
        "01111110" when "11110010",
        "00010000" when "11110011",
        "11000001" when "11110100",
        "10100101" when "11110101",
        "11001001" when "11110110",
        "00101111" when "11110111",
        "10010101" when "11111000",
        "11011000" when "11111001",
        "11000110" when "11111010",
        "10101100" when "11111011",
        "01100000" when "11111100",
        "01100100" when "11111101",
        "10101111" when "11111110",
        "00000000" when "11111111",
        "--------" when others;    
        
end architecture;
